entity bin2gray_v1 is
	port
	(
		b0, b1, b2, b3  : in bit;
		g0, g1, g2, g3  : in bit
	);
end entity;
--Exemplo implementando o circuito diretamente com as portas lógicas
architecture ifsc_v1 of bin2gray_v1 is
begin

end architecture;